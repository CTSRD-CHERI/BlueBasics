{-
 - Copyright (c) 2018-2019 Alexandre Joannou
 - All rights reserved.
 -
 - This software was developed by SRI International and the University of
 - Cambridge Computer Laboratory (Department of Computer Science and
 - Technology) under DARPA contract HR0011-18-C-0016 ("ECATS"), as part of the
 - DARPA SSITH research programme.
 -
 - @BERI_LICENSE_HEADER_START@
 -
 - Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 - license agreements.  See the NOTICE file distributed with this work for
 - additional information regarding copyright ownership.  BERI licenses this
 - file to you under the BERI Hardware-Software License, Version 1.0 (the
 - "License"); you may not use this file except in compliance with the
 - License.  You may obtain a copy of the License at:
 -
 -   http://www.beri-open-systems.org/legal/license-1-0.txt
 -
 - Unless required by applicable law or agreed to in writing, Work distributed
 - under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 - CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 - specific language governing permissions and limitations under the License.
 -
 - @BERI_LICENSE_HEADER_END@
 -}

package MasterSlave where

import SourceSink
import Connectable

-------------------------------
-- Master / Slave interfaces --
--------------------------------------------------------------------------------

interface Master req resp =
  source :: Source req
  sink   :: Sink resp

interface Slave req resp =
  source :: Source resp
  sink   :: Sink req

---------------------------
-- Connectable instances --
--------------------------------------------------------------------------------

instance Connectable (Master req resp) (Slave req resp) where
  mkConnection m s = module mkConnection m.source s.sink
                            mkConnection s.source m.sink

instance Connectable (Slave req resp) (Master req resp) where
  mkConnection s m = module mkConnection m.source s.sink
                            mkConnection s.source m.sink

-----------
-- Utils --
--------------------------------------------------------------------------------
-- Get desired Master / Slave sub-interface
getMasterSource :: Master a b -> Source a
getMasterSource m = m.source
getMasterSink   :: Master a b -> Sink b
getMasterSink   m = m.sink
getSlaveSource  :: Slave a b -> Source b
getSlaveSource  s = s.source
getSlaveSink    :: Slave a b -> Sink a
getSlaveSink    s = s.sink
